-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: maria
-- 
-- Create Date:    01/06/2020 14:23:49
-- Project Name:   UControl
-- Module Name:    UControl.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity UControl is
	port(IR : in std_logic_vector(11 downto 0):= x"000";
	     senControl : out std_logic_vector(15 downto 0);
		 clk : in std_logic
		 );
end UControl;

architecture arq1 of UControl is

	type ROM is array (0 to 2047) of std_logic_vector(15 downto 0);
	constant Senales : ROM := (	x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 000
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 040
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 080-087   sum mem RF ----Suma
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 088
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 0A0-0A7
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 0A8-0AF   sum R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 0B0-0B7	sum R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 0B8-OBF	sum R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 0C0-0C7
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 0C8-0CF	sum R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 0D0-0D7	sum R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 0D8-0DF	sum R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 0E8-0EF	sum R1, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 0F0-0F7	sum R2, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 0F8-0FF	sum R3, #
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 100-107	Res mem, RF ----Resta
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 108-10F
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 110-117
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 118-11F
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 120-127
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 128-12F	Res R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 130-137	Res R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 138-13F	Res R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 140-147
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 148-14F   Res R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 150-157   Res R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 158-15F   Res R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 160-167
 								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 168-16F   Res R1,  #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 170-177   Res R2,  #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 178-17F   Res R3,  #
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 180-187   mul mem, RF ----Multiplicacion
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 188
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 190
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 198
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 1A0
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 1A8-1AF   mul R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 1B0-1B7   mul R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 1B8-1BF   mul R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 1C0                  0001 1100 0000
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 1C8-1CF   mul R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 1D0-1D7   mul R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 1D8-1DF   mul R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 1E0
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 1E8-1EF   mul R1,  #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 1F0-1F7   mul R2,  #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 1F8-1FF   mul R3,  #
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 200-207   div mem, RF ---- Division 
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 208
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 210
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 218
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 220
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 228-22F  div R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 230-237  div R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 238-23F  div R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 240
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 248-24F  div R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 250-257  div R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 258-25F  div R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 260
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 268-26F  div R1,  #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 270-277  div R2,  #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 278-27F  div R3,  #
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 280-287  AND mem, RF ----- AND
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 288
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 290
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 298
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 2A0
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 2A8-2AF  AND R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 2B0-2B7  AND R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 2B8-2BF  AND R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 2C0
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 2C8-2CF  AND R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 2D0-2D7  AND R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 2D8-2DF  AND R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 2E0
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 2E8-asd	AND R1, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 2F0
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 2F8
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 300-307	Or mem, RF				
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 308
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 310
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 318
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 320
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 328-32F`	Or R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 330-337	Or R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 338-33F	Or R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 340
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 348-34F	Or R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 350-357	Or R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 358-35F	Or R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 2E8-asd	OR R1, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 2F0
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 378-37F	Or R3, #	?
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 380
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 3A0
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 3A8-3AF	Not R1
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 3B0-3B7	Not R2
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 3B8-3BF	Not R3
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 3C0
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0120",x"00C0",  --- 400-407	Xor mem, RF		
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0009",x"0000",x"0000",x"0000",x"0000",  --- 428-42F	Xor R1, RF
								x"4000",x"2800",x"0400",x"0005",x"0000",x"0000",x"0000",x"0000",  --- 430-437	Xor R2, RF
								x"4000",x"2800",x"0400",x"0003",x"0000",x"0000",x"0000",x"0000",  --- 438-43F	Xor R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 440
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0009",x"0000",  --- 448-44F	Xor R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0005",x"0000",  --- 450-457	Xor R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0003",x"0000",  --- 458-45F	Xor R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0009",x"0000",  --- 2E8-asd	Xor R1, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0005",x"0000",  --- 2F0
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0003",x"0000",  --- 478-47F	Xor R3, #	?	
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 480
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0121",x"0060",  --- 500-507	Comp mem, RF					
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 508-50F
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0001",x"0000",x"0000",x"0000",x"0000",  --- 528-52F	Comp R1, RF
								x"4000",x"2800",x"0400",x"0001",x"0000",x"0000",x"0000",x"0000",  --- 530-537	Comp R2, RF
								x"4000",x"2800",x"0400",x"0001",x"0000",x"0000",x"0000",x"0000",  --- 538-53F	Comp R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 540
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0001",x"0000",  --- 548-54F	Comp R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0001",x"0000",  --- 550-557	Comp R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0001",x"0000",  --- 558-55F	Comp R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 560
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0001",x"0000",  --- 568-56F	Comp R1, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0001",x"0000",  --- 570-577	Comp R2, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0001",x"0000",  --- 578-57F	Comp R3, #
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0120",x"0060",x"0000",  --- 580-587	Move mem, RF			
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0008",x"0000",x"0000",x"0000",x"0000",  --- 5A8-5AF	Move R1, RF
								x"4000",x"2800",x"0400",x"0004",x"0000",x"0000",x"0000",x"0000",  --- 5B0-5B7	Move R2, RF
								x"4000",x"2800",x"0400",x"0002",x"0000",x"0000",x"0000",x"0000",  --- 5B8-5BF	Move R3, RF
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 5C0
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0008",x"0000",  --- 5C8-5CF	Move R1, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0004",x"0000",  --- 5D0-5D7	Move R2, mem
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0100",x"0002",x"0000",  --- 5D8-5DF	Move R3, mem
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0008",x"0000",  --- 5E8-5EF	Move R1, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0004",x"0000",  --- 5F0-5F7	Move R2, #
								x"4000",x"2800",x"0400",x"4000",x"2800",x"0110",x"0002",x"0000",  --- 5F8-5FF	Move R3, #
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 600	Read RD, Puerto
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0130",x"0008",x"0000",  --- 608	Read R1, Puerto
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0130",x"0004",x"0000",  --- 610	Read R2, Puerto
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0130",x"0002",x"0000",  --- 618	Read R3, Puerto
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0120",x"00C0",x"0000",  --- 640	
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0120",x"00C0",x"0000",  --- 648	Write Puerto, RD
								x"4000",x"2800",x"0400",x"4000",x"2200",x"0120",x"00C0",x"0000",   	
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  	
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",  --- 680	Jump dir
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 0C0
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",  --- 700	CJmpG			
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",  --- 720	CjmpE
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"4000",x"2800",x"1000",x"0000",x"0000",  --- 740	CjmpL
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 180	Halt
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 1C0 0001 1100 0000
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"4000",x"2800",x"0400",x"0000",x"0000",x"0000",x"0000",x"0000" );
	signal LinDir : integer range 0 to 2047 := 0;
	signal contador : std_logic_vector(2 downto 0):= "000";	 
	signal Direccion : std_logic_vector(10 downto 0):= "00000000000";	

begin

process(clk)
	Variable cuentaP : unsigned(2 downto 0):="000";
begin 
	if clk'event and clk ='1' then
		cuentaP := cuentaP + 1;
	end if;
	contador <= std_logic_vector(cuentaP);
end process;

Direccion <= IR(11 downto 4) & contador;
LinDir <= to_integer(unsigned(Direccion));
senControl <= Senales(LinDir);

end arq1;
