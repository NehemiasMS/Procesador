-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: Marian Meza
-- 
-- Create Date:    17/04/2020 11:07:33
-- Project Name:   ROM_programa
-- Module Name:    ROM_programa.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity ROM_programa is
   port(A: in std_logic_vector(8 downto 0);
		D: out std_logic_vector(11 downto 0)
		);
end ROM_programa;

architecture arq1 of ROM_programa is
	type ROM is array(0 to 511) of std_logic_vector(11 downto 0);
--	constant Programa : ROM := (x"BD0",x"00A",x"BE0",x"014",x"BF0",x"01E",x"104",x"000",  --- 000   ---- EL PROGRAMA
--								x"158",x"190",x"000",x"1D0",x"001",x"208",x"001",x"26C",
--								x"000",x"2A0",x"001",x"2E0",x"002",x"30C",x"002",x"374",
--								x"3B0",x"002",x"3F0",x"003",x"404",x"003",x"474",x"490",
--								x"003",x"4D0",x"002",x"508",x"000",x"56C",x"5A0",x"002",
--								x"5E0",x"00A",x"60C",x"001",x"674",x"6B0",x"002",x"6F0",
--								x"006",x"760",x"804",x"002",x"86C",x"8A0",x"002",x"8D0",
--								x"007",x"A08",x"003",x"A74",x"AB0",x"003",x"AEF",x"EE9",
--								x"B0C",x"000",x"B58",x"BA0",x"001",x"BF0",x"009",x"C20",  --- 040
--								x"000",x"C88",x"010",x"000",x"000",x"000",x"000",x"000",

	constant Programa : ROM := (x"BD0",x"000",x"BE0",x"020",x"1D0",x"010",x"A58",x"E80",  --- 000  ---- JUUUUMPS
								x"011",x"A58",x"E40",x"004",x"A58",x"E00",x"004",x"1D0",
								x"010",x"BD0",x"000",x"000",x"000",x"000",x"000",x"000",

--	constant Programa : ROM := (x"BD0",x"000",x"C90",x"010",x"BE0",x"001",x"CA0",x"010",  --- 000  ---- FIBONACCIIII
--								x"BF0",x"002",x"158",x"C84",x"010",x"164",x"C88",x"010",
--								x"1F0",x"002",x"AF0",x"00A",x"E00",x"00A",x"D00",x"016",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 040
								
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 080
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 0C0
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 100
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 140
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 180
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",  --- 1C0
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000",
								x"000",x"000",x"000",x"000",x"000",x"000",x"000",x"000");				
begin
	D <= Programa(to_integer(unsigned(A)));
end arq1;
