-------------------------------------------------------------------------------
--
-- Company : Universidad Miguel Hernandez
-- Engineer: maria
-- 
-- Create Date:    01/06/2020 12:06:03
-- Project Name:   RAM
-- Module Name:    RAM.vhd
-- Description:
--
-- Additional Comments:
--
-------------------------------------------------------------------------------

library IEEE;
use IEEE.std_logic_1164.all;  -- Para std_logic
use IEEE.numeric_std.all;     -- Para unsigned

entity RAM is
   port(Direccion : in std_logic_vector(8 downto 0):= "000000000";
--      Palabra: inout std_logic_vector(15 downto 0):= x"0000";
		DatosE : in std_logic_vector(15 downto 0):= x"0000";
		DatosS : out std_logic_vector(15 downto 0):= x"0000";
        RW, IOM: in std_logic);
end RAM;

architecture arq1 of RAM is
	type dRAM is array (0 to 511) of std_logic_vector(15 downto 0);
	signal contador : dRAM :=(	x"0002",x"0200",x"0100",x"030A",x"0000",x"0000",x"0000",x"0000",  --- 000
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 040
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 080
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 0C0
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 100
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 140
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 180
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",  --- 1C0
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",
								x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000",x"0000");
	signal LinDir : integer range 0 to 511 := 0;
								
begin

process(Direccion, DatosE, RW, LinDir)
begin

	LinDir <= to_integer(unsigned(Direccion));
	
	if IOM = '0' then
		if RW = '1' then
			contador(LinDir) <= DatosE;
		else 
			DatosS <= contador(LinDir);
		end if;
	else 
		DatosS <= "ZZZZZZZZZZZZZZZZ";
	end if;

end process;

end arq1;
